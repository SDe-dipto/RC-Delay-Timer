<Qucs Schematic 0.0.5>
<Properties>
  <View=0,0,800,800,1,0,0>
  <Grid=10,10,1>
  <DataSet=schmitt.dat>
  <DataDisplay=schmitt.dpl>
  <OpenDisplay=1>
</Properties>
<Symbol>
</Symbol>
<Components>
  <R R1 1 120 130 15 -26 0 1 "4.7k" 1 "26.85" 0 "european" 0>
  <R R2 1 300 130 -53 -26 0 3 "4.7k" 1 "26.85" 0 "european" 0>
  <GND * 1 120 280 0 0 0 0>
  <GND * 1 300 280 0 0 0 0>
  <R R3 1 250 180 -26 15 0 0 "47k" 1 "26.85" 0 "european" 0>
  <R R4 1 180 280 15 -26 0 1 "47k" 1 "26.85" 0 "european" 0>
  <GND * 1 180 370 0 0 0 0>
  <Vpulse Ve 1 180 340 18 -26 0 1 "-5 V" 1 "+5 V" 1 "0" 1 "210 us" 1 "100 us" 0 "100 us" 0>
  <_BJT T2 1 120 250 -64 -26 1 2 "npn" 1 "1e-16" 0 "1" 0 "1" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "1.5" 0 "0" 0 "2" 0 "100" 0 "1" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0.75" 0 "0.33" 0 "1p" 1 "0.75" 0 "0.33" 0 "1.0" 0 "0" 0 "0.75" 0 "0" 0 "0.5" 0 "0.1n" 1 "0.0" 0 "0.0" 0 "0.0" 0 "0.0" 0 "26.85" 0 "0.0" 0 "1.0" 0 "1.0" 0 "0.0" 0 "1.0" 0 "1.0" 0 "0.0" 0>
  <_BJT T3 1 300 250 8 -26 0 0 "npn" 1 "1e-16" 0 "1" 0 "1" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "1.5" 0 "0" 0 "2" 0 "100" 0 "1" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0" 0 "0.75" 0 "0.33" 0 "1p" 1 "0.75" 0 "0.33" 0 "1.0" 0 "0" 0 "0.75" 0 "0" 0 "0.5" 0 "0.1n" 1 "0.0" 0 "0.0" 0 "0.0" 0 "0.0" 0 "26.85" 0 "0.0" 0 "1.0" 0 "1.0" 0 "0.0" 0 "1.0" 0 "1.0" 0 "0.0" 0>
  <.TR TR1 1 400 220 0 51 0 0 "lin" 1 "0 us" 1 "210 us" 1 "100" 0 "Trapezoidal" 0 "2" 0 "1 ns" 0 "1e-16" 0 "150" 0 "0.001" 0 "1 pA" 0 "1 uV" 0 "26.85" 0 "1e-3" 0 "1e-6" 0 "1" 0>
  <GND * 1 400 160 0 0 0 0>
  <Vdc Vdd 1 400 130 18 -26 0 1 "5 V" 1>
</Components>
<Wires>
  <300 80 300 100 "" 0 0 0>
  <120 80 120 100 "" 0 0 0>
  <120 80 300 80 "" 0 0 0>
  <300 160 300 180 "" 0 0 0>
  <280 180 300 180 "" 0 0 0>
  <120 160 120 180 "" 0 0 0>
  <120 180 120 220 "" 0 0 0>
  <300 180 300 220 "" 0 0 0>
  <180 180 220 180 "" 0 0 0>
  <150 250 180 250 "" 0 0 0>
  <180 180 180 250 "" 0 0 0>
  <120 180 160 180 "" 0 0 0>
  <160 230 240 230 "" 0 0 0>
  <160 180 160 230 "" 0 0 0>
  <240 250 270 250 "" 0 0 0>
  <240 230 240 250 "" 0 0 0>
  <400 80 400 100 "" 0 0 0>
  <300 80 400 80 "" 0 0 0>
  <180 310 180 310 "Input" 113 330 0>
  <300 180 300 180 "Output" 330 150 0>
</Wires>
<Diagrams>
</Diagrams>
<Paintings>
  <Text 60 40 16 #000000 0 "Schmitt-Trigger.">
  <Text 320 350 12 #000000 0 "This Schmitt-Trigger switches on at 1.7V and\nswitches off at approximately -2.7V.">
</Paintings>